
class my_driver extends uvm_driver#(my_sequence_item);
  `uvm_component_utils(my_driver)
  
   my_sequence_item seq_item;
   virtual intf my_vif;
  
  function new(string name = "my_driver", uvm_component parent = null);
  super.new(name, parent);
  endfunction
  
  function void build_phase(uvm_phase phase);
  super.build_phase(phase);

   if(!uvm_config_db#(virtual intf)::get(this, "", "my_vif", my_vif))
      `uvm_fatal(get_full_name(), "Error")
       
  endfunction

  task run_phase(uvm_phase phase);
  super.run_phase(phase);

    forever begin
      seq_item_port.get_next_item(seq_item);

      @(negedge my_vif.clk);
  
      my_vif.cipher_key <= seq_item.cipher_key; 
      my_vif.plain_text <= seq_item.plain_text;
      my_vif.valid_in   <= seq_item.valid_in;
      my_vif.reset      <= seq_item.reset;

      seq_item_port.item_done();
    
    end
  endtask
  
endclass
